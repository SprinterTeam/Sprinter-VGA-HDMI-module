-- megafunction wizard: %ALTLVDS%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altlvds_tx 

-- ============================================================
-- File Name: serializer.vhd
-- Megafunction Name(s):
-- 			altlvds_tx
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.0 Build 235 06/17/2009 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY serializer IS
	PORT
	(
		tx_in		: IN STD_LOGIC_VECTOR (29 DOWNTO 0);
		tx_inclock		: IN STD_LOGIC  := '0';
		tx_syncclock		: IN STD_LOGIC  := '0';
		tx_out		: OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END serializer;


ARCHITECTURE SYN OF serializer IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (2 DOWNTO 0);



	COMPONENT altlvds_tx
	GENERIC (
		deserialization_factor		: NATURAL;
		implement_in_les		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		number_of_channels		: NATURAL;
		registered_input		: STRING;
		use_external_pll		: STRING
	);
	PORT (
			tx_out	: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			tx_in	: IN STD_LOGIC_VECTOR (29 DOWNTO 0);
			tx_syncclock	: IN STD_LOGIC ;
			tx_inclock	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	tx_out    <= sub_wire0(2 DOWNTO 0);

	altlvds_tx_component : altlvds_tx
	GENERIC MAP (
		deserialization_factor => 10,
		implement_in_les => "ON",
		intended_device_family => "Cyclone",
		lpm_type => "altlvds_tx",
		number_of_channels => 3,
		registered_input => "OFF",
		use_external_pll => "ON"
	)
	PORT MAP (
		tx_in => tx_in,
		tx_syncclock => tx_syncclock,
		tx_inclock => tx_inclock,
		tx_out => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: Deser_Factor NUMERIC "10"
-- Retrieval info: PRIVATE: Enable_DPA_Mode STRING "OFF"
-- Retrieval info: PRIVATE: Ext_PLL STRING "ON"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone"
-- Retrieval info: PRIVATE: Int_Device STRING "Cyclone"
-- Retrieval info: PRIVATE: LVDS_Mode NUMERIC "0"
-- Retrieval info: PRIVATE: Le_Serdes STRING "ON"
-- Retrieval info: PRIVATE: Num_Channel NUMERIC "3"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "10"
-- Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "ON"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_tx"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "3"
-- Retrieval info: CONSTANT: REGISTERED_INPUT STRING "OFF"
-- Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "ON"
-- Retrieval info: USED_PORT: tx_in 0 0 30 0 INPUT NODEFVAL tx_in[29..0]
-- Retrieval info: USED_PORT: tx_inclock 0 0 0 0 INPUT_CLK_EXT GND tx_inclock
-- Retrieval info: USED_PORT: tx_out 0 0 3 0 OUTPUT NODEFVAL tx_out[2..0]
-- Retrieval info: USED_PORT: tx_syncclock 0 0 0 0 INPUT GND tx_syncclock
-- Retrieval info: CONNECT: @tx_in 0 0 30 0 tx_in 0 0 30 0
-- Retrieval info: CONNECT: tx_out 0 0 3 0 @tx_out 0 0 3 0
-- Retrieval info: CONNECT: @tx_syncclock 0 0 0 0 tx_syncclock 0 0 0 0
-- Retrieval info: CONNECT: @tx_inclock 0 0 0 0 tx_inclock 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL serializer.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL serializer.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL serializer.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL serializer.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL serializer.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL serializer_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
